class calc_sb #(int DataSize, int AddrSize);

  // Signals needed for the golden model implementation in the scoreboard
  int mem_a [2**AddrSize];
  int mem_b [2**AddrSize];
  logic second_read = 0;
  int golden_lower_data;
  int golden_upper_data;
  mailbox #(calc_seq_item #(DataSize, AddrSize)) sb_box;

  function new(mailbox #(calc_seq_item #(DataSize, AddrSize)) sb_box);
    this.sb_box = sb_box;
  endfunction

  task main();
    calc_seq_item #(DataSize, AddrSize) trans;
    forever begin
      sb_box.get(trans);
      //Initialize the SRAMs in the scoreboard's local memory
      if (trans.initialize) begin
        if (trans.lower_data !== 'x) begin
          mem_a[trans.curr_rd_addr] = trans.lower_data;
        end
        if (trans.upper_data !== 'x) begin
          mem_b[trans.curr_rd_addr] = trans.upper_data;
        end
        $display($stime, " SB: Init SRAM B addr=0x%0x data=0x%0x", trans.curr_wr_addr, trans.upper_data);
      end
      continue;	
      end

    // Read Operations
    if (trans.rdn_wr == 0) begin
      if (!second_read) begin
        golden_lower_data = trans.lower_data;
        golden_upper_data = trans.upper_data;
        second_read = 1;
      end
      if (second_read) begin
        if ((

      // The scoreboard's task is to verify the DUT's behavior by comparing the
      // data received from the monitor against a golden reference model.

      // Use the transaction flags (`initialize`, `rdn_wr`) to handle three distinct operations:
      // - For initialization, update the scoreboard's local memory (`mem_a` and `mem_b`) to match the DUT's initial SRAM state.
      // - For read operations, ompare the data from the SRAM in the DUT to the data stored in the scoreboard's memory.
      //       Think about how to account for the two sequential reads in the DUT for the single write operation. The values
      //       from both read operations need to be used to compare against the calculated values in the DUT when they are written
      //       to SRAM. The second_read, golden_lower_data, and golden_upper_data signals can be used for this purpose.
      // - For write operations, compare the DUT's output to the data calculated by the golden model in the scoreboard.

      // Use `$display` to log successful transactions and `$error` to report mismatches.
      // If a mismatch occurs, use `$finish` to terminate the simulation.
    end
  endtask

endclass : calc_sb
